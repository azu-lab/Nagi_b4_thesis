import(<kernel.cdl>);

typedef int_t   pup_direction_t;
typedef int_t   pbio_port_id_t;
typedef int_t   pbio_error_t;
typedef int_t   pup_motor_t;
typedef int_t   pup_device_t;
typedef int_t   bool;

signature sMotor {
    void set_motor_ref( void );
    void setup( [in] pup_direction_t positive_direction, [in] bool reset_count );
    void set_speed( [in] int32_t speed );
    void stop( void );
};

signature sSensor {
    void set_device_ref( void );
    void get_distance( [out] int32_t* distance );
    void light_on( void );
    void light_set( [in] int32_t bv1, [in] int32_t bv2, [in] int32_t bv3, [in] int32_t bv4 );
    void light_off( void );
};

signature sPowerdown{
    void powerdown( [in] pbio_error_t error );
};

celltype tMotor {
    call sPowerdown cPowerdown;
    entry sMotor eMotor;
    attr {
        pbio_port_id_t port = C_EXP("PBIO_PORT_ID_$port$");
    };
    var {
       pup_motor_t *motor = C_EXP("NULL");
    };
};

celltype tSensor {
    call sPowerdown cPowerdown;
    entry sSensor eSensor;
    attr{
        pbio_port_id_t port = C_EXP("PBIO_PORT_ID_$port$");
    };
    var {
        pup_device_t ult = C_EXP("NULL");
    };
};

celltype tTaskbody {
    entry sTaskBody eTaskbody;
    call sSensor cSensor;
    call sMotor cMotor;
};

celltype tPowerdown {
    entry sPowerdown ePowerdown1;
    entry sPowerdown ePowerdown2;
};

cell tMotor Motor {
    cPowerdown = Powerdown.ePowerdown1;
    port = C_EXP("PBIO_PORT_ID_A");
};

cell tSensor Sensor {
    cPowerdown = Powerdown.ePowerdown2;
    port = C_EXP("PBIO_PORT_ID_B");
};

cell tTaskbody Taskbody {
    cMotor = Motor.eMotor;
    cSensor = Sensor.eSensor;
};

cell tPowerdown Powerdown{
};

cell tTask Task{
    cTaskBody = Taskbody.eTaskbody;
    id = C_EXP("TASK1");
    attribute = C_EXP("TA_ACT");
    stackSize = C_EXP("STACK_SIZE");
    priority = C_EXP("HIGH_PRIORITY");
};