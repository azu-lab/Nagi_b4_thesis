
/* typedef int32_t ER; */

signature sMain {
	void  main(void);
};

signature sSig1 {
	ER func1( [in]int32_t arg1, [out]int32_t *res );
};

signature sSig2 {
	ER func1( [in]int32_t arg1, [out]int32_t *res );
};

signature sSig3 {
	ER func1( [in]int32_t arg1, [out]int32_t *res );
};

celltype tCtR1 {
	entry sSig3 eEnt;
};

celltype tCtR2 {
	call sSig2 cCall2;
	call sSig3 cCall3;
	entry sSig1 eEnt;
};

celltype tCtOuter {
	call    sSig1  cCall;
	entry   sSig2  eEnt;
	entry   sMain  eMain;
};

// TracePlugin で使われる
cell tSysLog  SysLogn2{
};
cell tKernel  Kernel{
};

/* rRegion2 初出現で specifier を指定 */
[to_through(rRegion1),
//[to_through(rRegion1, TracePlugin, "cellEntry=\"r1cell.eEnt2 , r1cell.eEnt\""),
//[to_through(rRegion1, TracePlugin, "cellEntry=\"r1cell.eEnt2\",cellEntry=\"r1cell.eEnt\""),
//[to_through(rRegion1, TracePlugin, "cellEntry=\"r1cell.eEnt2\""),
out_through(/*TracePlugin,""*/),
in_through()]
region rRegion2 {
};

region rRegion2 {
	/* プロトタイプ宣言 */
	cell tCtR2 r2cell;
};

/* rRegion1 初出現で specifier を指定 */
[from_through(rRegion2, TracePlugin, ""), out_through()]
region rRegion1{
	/* プロトタイプ宣言 */
	cell tCtR1 r1cell;

	// TracePlugin で使われる
//	cell tSysLog  SysLogn1{
//	};
};

cell tCtOuter outer {
	cCall = rRegion2::r2cell.eEnt;
};

/* ここ（再出現）では specifier を指定できない */
region rRegion1 {
	cell tCtR1 r1cell {
	};
};

/* ここ（再出現）では specifier を指定できない */
region rRegion2 {
	cell tCtR2 r2cell {
		cCall2 = outer.eEnt;
		cCall3 = rRegion1::r1cell.eEnt;
	};

	[out_through(Plugin2,"")]
	region rRegionInner {
		cell tCtR2 r2cellInner {
			cCall2 = outer.eEnt;
			/* #327 呼び口の through が region の through よりも前に出ることのテスト */
			[through(Plugin1, "" )]
				cCall3 = rRegion1::r1cell.eEnt;
		};
	};
};

[singleton,active]
celltype tMain {
	call sMain cMain;
};

cell tMain Main{
	cMain = outer.eMain;
};

