//import( <cygwin_kernel.cdl> );

//[deviate]
//signature sAllocator {
//   void  alloc( [in]int32_t size, [out]void **buf );
//   void  dealloc( [in]const void *buf );
//};

//celltype tAllocator {
//    entry  sAllocator eAlloc;
//};

//cell tAllocator Allocator {};

//cell tAllocator Allocator2 {};


//[generate( RustGenPlugin, "")]
signature sSample {
    void  print ( [in]int8_t varin, [out]int32_t *varout, [out]int32_t *varout2);
};

signature sSample2 {
	void print ([in,string(256)]const char_t *buf_in, [out,string(len)]char_t *buf_out, [in]int32_t len );
};

[generate( RustGenPlugin, "")]
celltype tSample {
	call sSample cPrint;
	call sSample2 cPrint2;
//	call sSample cPrint2;
};

[generate( RustGenPlugin, "")]
celltype tPrint {
	entry sSample ePrint;
	entry sSample2 ePrint2;
	call sSample cCalculate;
	attr{
        int16_t attribute = 1;
    };
    var {
		int16_t variable = 0;
	};
};

[generate(RustGenPlugin, "")]
celltype tCalculate {
	entry sSample eCalculate;
	attr{
		int32_t attribute = 4;
	};
	var{
		int32_t variable = 3;
	};
};

cell tCalculate Calcu{
};

//[generate( RustGenPlugin, "")]
//[allocator(ePrint.print.varsend=Allocator.eAlloc)]
cell tPrint PrintA {
	cCalculate = Calcu.eCalculate;
};

//[generate( RustGenPlugin, "")]
//cell tPrint PrintB {
//};

//[generate( RustGenPlugin, "")]
cell tSample Sample {
	cPrint = PrintA.ePrint;
	cPrint2 = PrintA.ePrint2;
//	cPrint2 = PrintB.ePrint;
};
