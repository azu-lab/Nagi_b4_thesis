// import(<kernel.cdl>);
import(<kernel_rs.cdl>);

[generate( RustGenPlugin, "")]
celltype tPrint {
	entry sTaskBody ePrint;
	call sTask cTask;
	attr{
		int32_t printattr = 1;
	};
	var{
		int32_t printvar = 10;
	};
};

[generate( RustGenPlugin, "")]
cell tPrint PrintA{
	cTask = Task.eTask;
	printattr = 2;
};

[generate( RustGenPlugin, "")]
cell tTask Task{
    cTaskBody = PrintA.ePrint;

    id = C_EXP("TASK1");
	//task = C_EXP("TASK1_REF");
	task_ref = C_EXP("unsafe{TaskRef::from_raw_nonnull(NonZeroI32::new(TASK1).unwrap())}");
    attribute = C_EXP("TA_ACT");
    stackSize = 1024;
    priority = 42;
};

