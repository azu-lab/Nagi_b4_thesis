import(<kernel_rs.cdl>);

typedef int_t   bool;

signature sBinarySearch {
	int32_t binary_search( [in] int32_t key);
};

signature sCompare {
	void cmp( [in] int32_t value, [in] int32_t key, [out] int32_t *left, [out] int32_t *right, [in] int32_t mind );
};

[generate( RustGenPlugin, "lib")]
celltype tTaskBody {
	entry sTaskBody eTaskbody;
	call sBinarySearch cBinarySearch;
	attr {
		int32_t key = 0;
	};
};

[generate( RustGenPlugin, "lib")]
celltype tBinarySearch {
	entry sBinarySearch eBinarySearch;
	call sCompare cCompare;
	attr {
        [size_is(100)]
            int32_t *array = {1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100};
	};
	var {
		int32_t left = 0;
		int32_t right = 99;
	};
};

[generate( RustGenPlugin, "lib")]
celltype tCompare {
	entry sCompare eCompare;
};

cell tTaskBody Taskbody {
	cBinarySearch = Binarysearch.eBinarySearch;
	key = 77;
};

cell tBinarySearch Binarysearch {
	cCompare = Compare.eCompare;
};

cell tCompare Compare {
};

[generate( ItronrsGenPlugin, "lib")]
cell tTask_rs Task{
    cTaskBody = Taskbody.eTaskbody;
    id = C_EXP("TASK1");
	task_ref = C_EXP("unsafe{TaskRef::from_raw_nonnull(NonZeroI32::new(TASK1).unwrap())}");
    attribute = C_EXP("TA_ACT");
    stackSize = 1024;
    priority = 42;
};